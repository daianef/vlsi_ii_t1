///////////////////////////////////////////////////////////////////////////////
// Copyright 2003 DEIS - Universita' di Bologna
// 
// name         testbenchtlm.v
// author       Federico Angiolini - fangiolini@deis.unibo.it
// info         Script to achieve xpipes platform synthesis.
//
///////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////
//           Automatically generated by xpipesCompiler - don't edit          //
//                File generated for topology: switch6x4power                //
///////////////////////////////////////////////////////////////////////////////

`timescale 1 ns / 1 ns
`include "settings.v"
`include "./switch_power_defines.v"

module testbench();
  
  // May be overridden by the simulation scripts
  parameter TESTINGMODE = `ROTATE;
  parameter FLITWIDTH = 67;
  parameter NUMBERINPUTS = 6;
  parameter LOGNUMBERINPUTS = 3;
  parameter NUMBEROUTPUTS = 6;
  parameter LOGNUMBEROUTPUTS = 3;
  parameter CLOCKSEMIPERIOD = 2500;
  // The SIMDELAY knob is used at the interface between behavioural-style traffic generators and netlist-level representation of the topology under
  // test. The delay should be set so as to respect setup/propagation times at the input/output pins of the netlist, and be shorter than the clock period.
  parameter SIMDELAY = CLOCKSEMIPERIOD * 0.4;
  
  reg                           clk;
  reg                           rst;
  reg [LOGNUMBERINPUTS - 1:0]   ID [NUMBERINPUTS - 1:0];
  
  wire [FLITWIDTH - 1:0]        FLIT_in [NUMBERINPUTS - 1:0];
  wire                          VALID_in [NUMBERINPUTS - 1:0];
  wire                          FWDAUX1_in [NUMBERINPUTS - 1:0];
  wire                          BWDAUX1_out [NUMBERINPUTS - 1:0];
  wire                          BWDAUX2_out [NUMBERINPUTS - 1:0];
  wire                          BWDAUX3_out [NUMBERINPUTS - 1:0];
  
  wire [FLITWIDTH - 1:0]        FLIT_out [NUMBEROUTPUTS - 1:0];
  wire                          VALID_out [NUMBEROUTPUTS - 1:0];
  wire                          FWDAUX1_out [NUMBEROUTPUTS - 1:0];
  wire                          BWDAUX1_in [NUMBEROUTPUTS - 1:0];
  wire                          BWDAUX2_in [NUMBEROUTPUTS - 1:0];
  wire                          BWDAUX3_in [NUMBEROUTPUTS - 1:0];
  
  integer                       loop;
  
  genvar                        i;
  
  generate
    begin
      for (i = 0; i < NUMBERINPUTS; i = i + 1)
        begin : tester_input
          switch_power_tester_input #(.TESTINGMODE(TESTINGMODE), .FLITWIDTH(FLITWIDTH), .NUMBERINPUTS(NUMBERINPUTS), .LOGNUMBERINPUTS(LOGNUMBERINPUTS), .NUMBEROUTPUTS(NUMBEROUTPUTS), .LOGNUMBEROUTPUTS(LOGNUMBEROUTPUTS), .SIMDELAY(SIMDELAY))
                                    ti(clk, rst, ID[i],
                                       FLIT_in[i], VALID_in[i], FWDAUX1_in[i],
                                       BWDAUX1_out[i], BWDAUX2_out[i], BWDAUX3_out[i]);
        end
    end
  endgenerate
  
  generate
    begin
      for (i = 0; i < NUMBEROUTPUTS; i = i + 1)
        begin : tester_output
          switch_power_tester_output #(.TESTINGMODE(TESTINGMODE), .FLITWIDTH(FLITWIDTH), .SIMDELAY(SIMDELAY))
                                     to(clk, rst,
                                        FLIT_out[i], VALID_out[i], FWDAUX1_out[i],
                                        BWDAUX1_in[i], BWDAUX2_in[i], BWDAUX3_in[i]);
        end
    end
  endgenerate
  
switch_6x6_2_6 dut(.clk(clk), .rst(rst),
                .FLIT_in__0(FLIT_in[0]), .VALID_in__0(VALID_in[0]), .FWDAUX1_in__0(FWDAUX1_in[0]), 
		.BWDAUX1_out__0(BWDAUX1_out[0]), .BWDAUX2_out__0(BWDAUX2_out[0]), .BWDAUX3_out__0(BWDAUX3_out[0]),
                .FLIT_in__1(FLIT_in[1]), .VALID_in__1(VALID_in[1]), .FWDAUX1_in__1(FWDAUX1_in[1]), 
		.BWDAUX1_out__1(BWDAUX1_out[1]), .BWDAUX2_out__1(BWDAUX2_out[1]), .BWDAUX3_out__1(BWDAUX3_out[1]),
                .FLIT_in__2(FLIT_in[2]), .VALID_in__2(VALID_in[2]), .FWDAUX1_in__2(FWDAUX1_in[2]), 
		.BWDAUX1_out__2(BWDAUX1_out[2]), .BWDAUX2_out__2(BWDAUX2_out[2]), .BWDAUX3_out__2(BWDAUX3_out[2]),
                .FLIT_in__3(FLIT_in[3]), .VALID_in__3(VALID_in[3]), .FWDAUX1_in__3(FWDAUX1_in[3]), 
		.BWDAUX1_out__3(BWDAUX1_out[3]), .BWDAUX2_out__3(BWDAUX2_out[3]), .BWDAUX3_out__3(BWDAUX3_out[3]),
                .FLIT_in__4(FLIT_in[4]), .VALID_in__4(VALID_in[4]), .FWDAUX1_in__4(FWDAUX1_in[4]), 
		.BWDAUX1_out__4(BWDAUX1_out[4]), .BWDAUX2_out__4(BWDAUX2_out[4]), .BWDAUX3_out__4(BWDAUX3_out[4]),
                .FLIT_in__5(FLIT_in[5]), .VALID_in__5(VALID_in[5]), .FWDAUX1_in__5(FWDAUX1_in[5]), 
		.BWDAUX1_out__5(BWDAUX1_out[5]), .BWDAUX2_out__5(BWDAUX2_out[5]), .BWDAUX3_out__5(BWDAUX3_out[5]),
                .FLIT_out__0(FLIT_out[0]), .VALID_out__0(VALID_out[0]), .FWDAUX1_out__0(FWDAUX1_out[0]), 
		.BWDAUX1_in__0(BWDAUX1_in[0]), .BWDAUX2_in__0(BWDAUX2_in[0]), .BWDAUX3_in__0(BWDAUX3_in[0]),
                .FLIT_out__1(FLIT_out[1]), .VALID_out__1(VALID_out[1]), .FWDAUX1_out__1(FWDAUX1_out[1]), 
		.BWDAUX1_in__1(BWDAUX1_in[1]), .BWDAUX2_in__1(BWDAUX2_in[1]), .BWDAUX3_in__1(BWDAUX3_in[1]),
                .FLIT_out__2(FLIT_out[2]), .VALID_out__2(VALID_out[2]), .FWDAUX1_out__2(FWDAUX1_out[2]), 
		.BWDAUX1_in__2(BWDAUX1_in[2]), .BWDAUX2_in__2(BWDAUX2_in[2]), .BWDAUX3_in__2(BWDAUX3_in[2]),
                .FLIT_out__3(FLIT_out[3]), .VALID_out__3(VALID_out[3]), .FWDAUX1_out__3(FWDAUX1_out[3]), 
		.BWDAUX1_in__3(BWDAUX1_in[3]), .BWDAUX2_in__3(BWDAUX2_in[3]), .BWDAUX3_in__3(BWDAUX3_in[3]),
                .FLIT_out__4(FLIT_out[4]), .VALID_out__4(VALID_out[4]), .FWDAUX1_out__4(FWDAUX1_out[4]), 
		.BWDAUX1_in__4(BWDAUX1_in[4]), .BWDAUX2_in__4(BWDAUX2_in[4]), .BWDAUX3_in__4(BWDAUX3_in[4]),
                .FLIT_out__5(FLIT_out[5]), .VALID_out__5(VALID_out[5]), .FWDAUX1_out__5(FWDAUX1_out[5]), 
		.BWDAUX1_in__5(BWDAUX1_in[5]), .BWDAUX2_in__5(BWDAUX2_in[5]), .BWDAUX3_in__5(BWDAUX3_in[5]));
  
  
  initial
  begin
    // xpipes clock
    clk = 0;
    #(CLOCKSEMIPERIOD)
    forever #(CLOCKSEMIPERIOD) clk = ~clk;
  end
  

  initial
  begin
    // IDs
    for (loop = 0 ; loop < NUMBERINPUTS ; loop = 1 + loop)
      ID[loop] = loop;
  end
  
  initial
  begin
    rst = !`RESETACTIVEVALUE;
    #(2.5 * CLOCKSEMIPERIOD);
    rst = `RESETACTIVEVALUE;
    #(10 * CLOCKSEMIPERIOD);
    rst = !`RESETACTIVEVALUE;
  end
endmodule
